module ast

